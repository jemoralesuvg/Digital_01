module top();



endmodule
