
module top (
	input PIN_10, PIN_13, PIN_7,
	output PIN_14, PIN_17, PIN_20, PIN_23
);
	
	assign PIN_14 = PIN_10;
	
endmodule